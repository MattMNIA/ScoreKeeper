module	bcd_converter(N2,N1,X);
	input [4:0] X;
	output [3:0] N2;
	output [3:0] N1;
		assign N2[3] = 0;
		assign N2[2] = 0;
		assign N2[1] = (X[4]&X[3])|(X[4]&X[2]);
		assign N2[0] =((~X[4])&X[3]&X[1])|((~X[4])&X[3]&X[2])|(X[3]&X[2]&X[1])|(X[4]&(~X[3])&(~X[2])) ;
		assign N1[3] = ((~X[4])&X[3]&(~X[2])&(~X[1]))|(X[4]&(~X[3])&(~X[2])&X[1])|(X[4]&X[3]&X[2]&(~X[1]));
		assign N1[2] =((~X[4])&(~X[3])&X[2])|((~X[4])&X[2]&X[1])|(X[4]&(~X[2])&(~X[1]))|(X[4]&X[3]&(~X[2])) ;
		assign N1[1] = ((~X[4])&(~X[3])&(X[1]))|((~X[3])&X[2]&X[1])|((~X[4])&X[3]&X[2]&(~X[1]))|(X[4]&(~X[3])&(~X[2])&(~X[1]))|(X[4]&X[3]&(~X[2])&X[1]);
		assign N1[0] = X[0];
endmodule