module seven_seg_decoder(A, B, C, D, E, F, G, X);
	input [3:0] X;
	output A, B, C, D, E, F, G;
		assign A = (~X[3]&~X[2]&~X[1]&X[0])| (~X[3]&X[2]&~X[1]&~X[0])| (X[3]&X[2]&~X[1]&X[0])|(X[3]&~X[2]&X[1]&X[0]);
		assign B = (X[3]&X[1]&X[0])|(X[2]&X[1]&~X[0])|(X[3]&X[2]&~X[0])|(~X[3]&X[2]&~X[1]&X[0]);
		assign C = (X[3]&X[2]&X[1])|(X[3]&X[2]&~X[0])|(~X[3]&~X[2]&X[1]&~X[0]);
		assign D = (X[2]&X[1]&X[0])|(~X[3]&~X[2]&~X[1]&X[0])|( ~X[3]&X[2]&~X[1]&~X[0])|(X[3]&~X[2]&X[1]&~X[0]);
		assign E = (~X[3]&X[0])|(~X[2]&~X[1]&X[0])|(~X[3]&X[2]&~X[1]);
		assign F = (~X[3]&X[1]&X[0])|(~X[3]&~X[2]&X[0])|(~X[3]&~X[2]&X[1])|(X[3]&X[2]&~X[1]&X[0]);
		assign G = (~X[3]&~X[2]&~X[1])|(~X[3]&X[2]&X[1]&X[0])|( X[3]&X[2]&~X[1]&~X[0]);
endmodule